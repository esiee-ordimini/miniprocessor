library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity compteur_point is
port (
	-----------------------------------------------------------------
	-- Signaux d'affichage
	-----------------------------------------------------------------
	point_hexa 			: in std_logic_vector(9 downto 0 );
	point_dec			: out std_logic_vector(24 downto 0);

);
end entity;

architecture rtl of compteur_point is
begin

process(point_hexa)
 begin
  case point_hexa is
	when "000000000" => abcdefg <= "0000 0000 0000 0000 0000 0000";  -- 0
    when "000000001" => abcdefg <= "0000 0000 0000 0000 0000 0001";  -- 1
    when "000000010" => abcdefg <= "0000 0000 0000 0000 0000 0010";  -- 2
    when "000000011" => abcdefg <= "0000 0000 0000 0000 0000 0011";  -- 3
    when "000000100" => abcdefg <= "0000 0000 0000 0000 0000 0100";  -- 4
    when "000000101" => abcdefg <= "0000 0000 0000 0000 0000 0101";  -- 5
    when "000000110" => abcdefg <= "0000 0000 0000 0000 0000 0110";  -- 6
    when "000000111" => abcdefg <= "0000 0000 0000 0000 0000 0111";  -- 7
    when "000001000" => abcdefg <= "0000 0000 0000 0000 0000 1000";  -- 8
    when "000001001" => abcdefg <= "0000 0000 0000 0000 0000 1001";  -- 9
    when "000001010" => abcdefg <= "0000 0000 0000 0000 0001 0000";  -- 10
    when "000001011" => abcdefg <= "0000 0000 0000 0000 0001 0001";  -- 11
    when "000001100" => abcdefg <= "0000 0000 0000 0000 0001 0010";  -- 12
    when "000001101" => abcdefg <= "0000 0000 0000 0000 0001 0011";  -- 13
    when "000001110" => abcdefg <= "0000 0000 0000 0000 0001 0100";  -- 14
    when "000001111" => abcdefg <= "0000 0000 0000 0000 0001 0101";  -- 15
	when "000010001" => abcdefg <= "0000 0000 0000 0000 0001 0110";  -- 16
    when "000010010" => abcdefg <= "0000 0000 0000 0000 0001 0111";  -- 17
    when "000010011" => abcdefg <= "0000 0000 0000 0000 0001 1000";  -- 18
    when "000010100" => abcdefg <= "0000 0000 0000 0000 0001 1001";  -- 19
	 
	when "000010101" => abcdefg <= "0000 0000 0000 0000 0010 0000";  -- 20
    when "000010110" => abcdefg <= "0000 0000 0000 0000 0010 0001";  -- 21
    when "000010111" => abcdefg <= "0000 0000 0000 0000 0010 0010";  -- 22
    when "000011000" => abcdefg <= "0000 0000 0000 0000 0010 0011";  -- 23
    when "000011001" => abcdefg <= "0000 0000 0000 0000 0010 0100";  -- 24
    when "000011010" => abcdefg <= "0000 0000 0000 0000 0010 0101";  -- 25
    when "000011011" => abcdefg <= "0000 0000 0000 0000 0010 0110";  -- 26
    when "000011100" => abcdefg <= "0000 0000 0000 0000 0010 0111";  -- 27
    when "000011101" => abcdefg <= "0000 0000 0000 0000 0010 1000";  -- 28
    when "000011110" => abcdefg <= "0000 0000 0000 0000 0010 1001";  -- 29
    when "000011111" => abcdefg <= "0000 0000 0000 0000 0011 0000";  -- 30
    when "000100000" => abcdefg <= "0000 0000 0000 0000 0011 0001";  -- 31
    when "000100001" => abcdefg <= "0000 0000 0000 0000 0011 0010";  -- 32
    when "000100010" => abcdefg <= "0000 0000 0000 0000 0011 0011";  -- 33
    when "000100011" => abcdefg <= "0000 0000 0000 0000 0011 0100";  -- 34
    when "000100100" => abcdefg <= "0000 0000 0000 0000 0011 0101";  -- 35
	when "000100101" => abcdefg <= "0000 0000 0000 0000 0011 0110";  -- 36
    when "000100110" => abcdefg <= "0000 0000 0000 0000 0011 0111";  -- 37
    when "000100111" => abcdefg <= "0000 0000 0000 0000 0011 1000";  -- 38
    when "000101000" => abcdefg <= "0000 0000 0000 0000 0011 1001";  -- 39

	when "000101001" => abcdefg <= "0000 0000 0000 0000 0100 0000";  -- 40
    when "000101010" => abcdefg <= "0000 0000 0000 0000 0100 0001";  -- 41
    when "000101011" => abcdefg <= "0000 0000 0000 0000 0100 0010";  -- 42
    when "000101100" => abcdefg <= "0000 0000 0000 0000 0100 0011";  -- 43
    when "000101101" => abcdefg <= "0000 0000 0000 0000 0100 0100";  -- 44
    when "000101110" => abcdefg <= "0000 0000 0000 0000 0100 0101";  -- 45
    when "000101111" => abcdefg <= "0000 0000 0000 0000 0100 0110";  -- 46
    when "000110001" => abcdefg <= "0000 0000 0000 0000 0100 0111";  -- 47
    when "000110010" => abcdefg <= "0000 0000 0000 0000 0100 1000";  -- 48
    when "000110011" => abcdefg <= "0000 0000 0000 0000 0100 1001";  -- 49
    when "000110100" => abcdefg <= "0000 0000 0000 0000 0101 0000";  -- 50
    when "000110101" => abcdefg <= "0000 0000 0000 0000 0101 0001";  -- 51
    when "000110110" => abcdefg <= "0000 0000 0000 0000 0101 0010";  -- 52
    when "000110111" => abcdefg <= "0000 0000 0000 0000 0101 0011";  -- 53
    when "000111000" => abcdefg <= "0000 0000 0000 0000 0101 0100";  -- 54
    when "000111001" => abcdefg <= "0000 0000 0000 0000 0101 0101";  -- 55
	when "000111010" => abcdefg <= "0000 0000 0000 0000 0101 0110";  -- 56
    when "000111011" => abcdefg <= "0000 0000 0000 0000 0101 0111";  -- 57
    when "000111100" => abcdefg <= "0000 0000 0000 0000 0101 1000";  -- 58
    when "000111101" => abcdefg <= "0000 0000 0000 0000 0101 1001";  -- 59

	when "000111111" => abcdefg <= "0000 0000 0000 0000 0100 0000";  -- 60
    when "001000001" => abcdefg <= "0000 0000 0000 0000 0100 0001";  -- 61
    when "001000010" => abcdefg <= "0000 0000 0000 0000 0100 0010";  -- 62
    when "001000011" => abcdefg <= "0000 0000 0000 0000 0100 0011";  -- 63
    when "001000100" => abcdefg <= "0000 0000 0000 0000 0100 0100";  -- 64
    when "001000101" => abcdefg <= "0000 0000 0000 0000 0100 0101";  -- 65
    when "001000110" => abcdefg <= "0000 0000 0000 0000 0100 0110";  -- 66
    when "001000111" => abcdefg <= "0000 0000 0000 0000 0100 0111";  -- 67
    when "001001000" => abcdefg <= "0000 0000 0000 0000 0100 1000";  -- 68
    when "001001001" => abcdefg <= "0000 0000 0000 0000 0100 1001";  -- 69
    when "001001010" => abcdefg <= "0000 0000 0000 0000 0101 0000";  -- 70
    when "001001011" => abcdefg <= "0000 0000 0000 0000 0101 0001";  -- 71
    when "001001100" => abcdefg <= "0000 0000 0000 0000 0101 0010";  -- 72
    when "001001101" => abcdefg <= "0000 0000 0000 0000 0101 0011";  -- 73
    when "001001110" => abcdefg <= "0000 0000 0000 0000 0101 0100";  -- 74
    when "001001111" => abcdefg <= "0000 0000 0000 0000 0101 0101";  -- 75
	when "001010000" => abcdefg <= "0000 0000 0000 0000 0101 0110";  -- 76
    when "001010001" => abcdefg <= "0000 0000 0000 0000 0101 0111";  -- 77
    when "001010010" => abcdefg <= "0000 0000 0000 0000 0101 1000";  -- 78
    when "001010011" => abcdefg <= "0000 0000 0000 0000 0101 1001";  -- 79

	when "001010100" => abcdefg <= "0000 0000 0000 0000 0100 0000";  -- 80
    when "001010101" => abcdefg <= "0000 0000 0000 0000 0100 0001";  -- 81
    when "001010110" => abcdefg <= "0000 0000 0000 0000 0100 0010";  -- 82
    when "001010111" => abcdefg <= "0000 0000 0000 0000 0100 0011";  -- 83
    when "001011000" => abcdefg <= "0000 0000 0000 0000 0100 0100";  -- 84
    when "001011001" => abcdefg <= "0000 0000 0000 0000 0100 0101";  -- 85
    when "001011010" => abcdefg <= "0000 0000 0000 0000 0100 0110";  -- 86
    when "001011011" => abcdefg <= "0000 0000 0000 0000 0100 0111";  -- 87
    when "001011100" => abcdefg <= "0000 0000 0000 0000 0100 1000";  -- 88
    when "001011101" => abcdefg <= "0000 0000 0000 0000 0100 1001";  -- 89
    when "001011110" => abcdefg <= "0000 0000 0000 0000 0101 0000";  -- 90
    when "001011111" => abcdefg <= "0000 0000 0000 0000 0101 0001";  -- 91
    when "001100000" => abcdefg <= "0000 0000 0000 0000 0101 0010";  -- 92
    when "001100001" => abcdefg <= "0000 0000 0000 0000 0101 0011";  -- 93
    when "001100010" => abcdefg <= "0000 0000 0000 0000 0101 0100";  -- 94
    when "001100011" => abcdefg <= "0000 0000 0000 0000 0101 0101";  -- 95
	when "001100100" => abcdefg <= "0000 0000 0000 0000 0101 0110";  -- 96
    when "001100101" => abcdefg <= "0000 0000 0000 0000 0101 0111";  -- 97
    when "001100110" => abcdefg <= "0000 0000 0000 0000 0101 1000";  -- 98
    when "001100111" => abcdefg <= "0000 0000 0000 0000 0101 1001";  -- 99


  end case;
 end process;

	
end architecture;