library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity compteur_point is
port (
	-----------------------------------------------------------------
	-- Signaux d'affichage
	-----------------------------------------------------------------
	point_hexa 			: in std_logic_vector(6 downto 0 );
	point_dec			: out std_logic_vector(24 downto 0)

);
end entity;

architecture rtl of compteur_point is
	signal abcdefg 			: std_logic_vector(23 downto 0);
begin

process(point_hexa)
 begin
  case point_hexa is
    when "0000000" => abcdefg <= "000000000000000000000000";  -- 0
    when "0000001" => abcdefg <= "000000000000000000000001";  -- 1
    when "0000010" => abcdefg <= "000000000000000000000010";  -- 2
    when "0000011" => abcdefg <= "000000000000000000000011";  -- 3
    when "0000100" => abcdefg <= "000000000000000000000100";  -- 4
    when "0000101" => abcdefg <= "000000000000000000000101";  -- 5
    when "0000110" => abcdefg <= "000000000000000000000110";  -- 6
    when "0000111" => abcdefg <= "000000000000000000000111";  -- 7
    when "0001000" => abcdefg <= "000000000000000000001000";  -- 8
    when "0001001" => abcdefg <= "000000000000000000001001";  -- 9
    when "0001010" => abcdefg <= "000000000000000000010000";  -- 10
    when "0001011" => abcdefg <= "000000000000000000010001";  -- 11
    when "0001100" => abcdefg <= "000000000000000000010010";  -- 12
    when "0001101" => abcdefg <= "000000000000000000010011";  -- 13
    when "0001110" => abcdefg <= "000000000000000000010100";  -- 14
    when "0001111" => abcdefg <= "000000000000000000010101";  -- 15
    when "0010001" => abcdefg <= "000000000000000000010110";  -- 16
    when "0010010" => abcdefg <= "000000000000000000010111";  -- 17
    when "0010011" => abcdefg <= "000000000000000000011000";  -- 18
    when "0010100" => abcdefg <= "000000000000000000011001";  -- 19
	 
    when "0010101" => abcdefg <= "000000000000000000100000";  -- 20
    when "0010110" => abcdefg <= "000000000000000000100001";  -- 21
    when "0010111" => abcdefg <= "000000000000000000100010";  -- 22
    when "0011000" => abcdefg <= "000000000000000000100011";  -- 23
    when "0011001" => abcdefg <= "000000000000000000100100";  -- 24
    when "0011010" => abcdefg <= "000000000000000000100101";  -- 25
    when "0011011" => abcdefg <= "000000000000000000100110";  -- 26
    when "0011100" => abcdefg <= "000000000000000000100111";  -- 27
    when "0011101" => abcdefg <= "000000000000000000101000";  -- 28
    when "0011110" => abcdefg <= "000000000000000000101001";  -- 29
    when "0011111" => abcdefg <= "000000000000000000110000";  -- 30
    when "0100000" => abcdefg <= "000000000000000000110001";  -- 31
    when "0100001" => abcdefg <= "000000000000000000110010";  -- 32
    when "0100010" => abcdefg <= "000000000000000000110011";  -- 33
    when "0100011" => abcdefg <= "000000000000000000110100";  -- 34
    when "0100100" => abcdefg <= "000000000000000000110101";  -- 35
    when "0100101" => abcdefg <= "000000000000000000110110";  -- 36
    when "0100110" => abcdefg <= "000000000000000000110111";  -- 37
    when "0100111" => abcdefg <= "000000000000000000111000";  -- 38
    when "0101000" => abcdefg <= "000000000000000000111001";  -- 39

    when "0101001" => abcdefg <= "000000000000000001000000";  -- 40
    when "0101010" => abcdefg <= "000000000000000001000001";  -- 41
    when "0101011" => abcdefg <= "000000000000000001000010";  -- 42
    when "0101100" => abcdefg <= "000000000000000001000011";  -- 43
    when "0101101" => abcdefg <= "000000000000000001000100";  -- 44
    when "0101110" => abcdefg <= "000000000000000001000101";  -- 45
    when "0101111" => abcdefg <= "000000000000000001000110";  -- 46
    when "0110001" => abcdefg <= "000000000000000001000111";  -- 47
    when "0110010" => abcdefg <= "000000000000000001001000";  -- 48
    when "0110011" => abcdefg <= "000000000000000001001001";  -- 49
    when "0110100" => abcdefg <= "000000000000000001010000";  -- 50
    when "0110101" => abcdefg <= "000000000000000001010001";  -- 51
    when "0110110" => abcdefg <= "000000000000000001010010";  -- 52
    when "0110111" => abcdefg <= "000000000000000001010011";  -- 53
    when "0111000" => abcdefg <= "000000000000000001010100";  -- 54
    when "0111001" => abcdefg <= "000000000000000001010101";  -- 55
    when "0111010" => abcdefg <= "000000000000000001010110";  -- 56
    when "0111011" => abcdefg <= "000000000000000001010111";  -- 57
    when "0111100" => abcdefg <= "000000000000000001011000";  -- 58
    when "0111101" => abcdefg <= "000000000000000001011001";  -- 59

    when "0111111" => abcdefg <= "000000000000000001000000";  -- 60
    when "1000001" => abcdefg <= "000000000000000001000001";  -- 61
    when "1000010" => abcdefg <= "000000000000000001000010";  -- 62
    when "1000011" => abcdefg <= "000000000000000001000011";  -- 63
    when "1000100" => abcdefg <= "000000000000000001000100";  -- 64
    when "1000101" => abcdefg <= "000000000000000001000101";  -- 65
    when "1000110" => abcdefg <= "000000000000000001000110";  -- 66
    when "1000111" => abcdefg <= "000000000000000001000111";  -- 67
    when "1001000" => abcdefg <= "000000000000000001001000";  -- 68
    when "1001001" => abcdefg <= "000000000000000001001001";  -- 69
    when "1001010" => abcdefg <= "000000000000000001010000";  -- 70
    when "1001011" => abcdefg <= "000000000000000001010001";  -- 71
    when "1001100" => abcdefg <= "000000000000000001010010";  -- 72
    when "1001101" => abcdefg <= "000000000000000001010011";  -- 73
    when "1001110" => abcdefg <= "000000000000000001010100";  -- 74
    when "1001111" => abcdefg <= "000000000000000001010101";  -- 75
    when "1010000" => abcdefg <= "000000000000000001010110";  -- 76
    when "1010001" => abcdefg <= "000000000000000001010111";  -- 77
    when "1010010" => abcdefg <= "000000000000000001011000";  -- 78
    when "1010011" => abcdefg <= "000000000000000001011001";  -- 79

    when "1010100" => abcdefg <= "000000000000000001000000";  -- 80
    when "1010101" => abcdefg <= "000000000000000001000001";  -- 81
    when "1010110" => abcdefg <= "000000000000000001000010";  -- 82
    when "1010111" => abcdefg <= "000000000000000001000011";  -- 83
    when "1011000" => abcdefg <= "000000000000000001000100";  -- 84
    when "1011001" => abcdefg <= "000000000000000001000101";  -- 85
    when "1011010" => abcdefg <= "000000000000000001000110";  -- 86
    when "1011011" => abcdefg <= "000000000000000001000111";  -- 87
    when "1011100" => abcdefg <= "000000000000000001001000";  -- 88
    when "1011101" => abcdefg <= "000000000000000001001001";  -- 89
    when "1011110" => abcdefg <= "000000000000000001010000";  -- 90
    when "1011111" => abcdefg <= "000000000000000001010001";  -- 91
    when "1100000" => abcdefg <= "000000000000000001010010";  -- 92
    when "1100001" => abcdefg <= "000000000000000001010011";  -- 93
    when "1100010" => abcdefg <= "000000000000000001010100";  -- 94
    when "1100011" => abcdefg <= "000000000000000001010101";  -- 95
    when "1100100" => abcdefg <= "000000000000000001010110";  -- 96
    when "1100101" => abcdefg <= "000000000000000001010111";  -- 97
    when "1100110" => abcdefg <= "000000000000000001011000";  -- 98
    when "1100111" => abcdefg <= "000000000000000001011001";  -- 99
    when others => abcdefg <= "111111111111111111111111";

  end case;
 end process;

	
end architecture;